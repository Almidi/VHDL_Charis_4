--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   18:12:26 02/12/2017
-- Design Name:   
-- Module Name:   C:/Users/JARVIS/Dropbox/ORGANWSH/Lab1/B/RF/DecoderUnitTest.vhd
-- Project Name:  RF
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: Decoder5x32
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY DecoderUnitTest IS
END DecoderUnitTest;
 
ARCHITECTURE behavior OF DecoderUnitTest IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT Decoder5x32
    PORT(
         Input : IN  std_logic_vector(4 downto 0);
         Output : OUT  std_logic_vector(31 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal Input : std_logic_vector(4 downto 0) := (others => '0');

 	--Outputs
   signal Output : std_logic_vector(31 downto 0);
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
   
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: Decoder5x32 PORT MAP (
          Input => Input,
          Output => Output
        );

   
 

    -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	
		Input<="00000";
		
		wait for 100 ns;
		Input<="00001";
		
		wait for 100 ns;
		Input<="00010";
		
		wait for 100 ns;

      -- insert stimulus here 

      wait;
   end process;

END;
